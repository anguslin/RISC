module decoder(instruction, nsel, opcode, readnum, writenum, ALUop, op, shift, sximm5, sximm8);
        //inputs and outputs
        input[15:0] instruction;
        input [2:0] nsel;
        output [2:0] opcode, readnum, writenum;
        output [1:0] ALUop, op, shift;
        output [15:0] sximm5, sximm8;

module datapath(clk, readnum, vsel, loada, loadb, shift, asel, bsel, ALUop, loadc, loads, writenum, write, mdata, sximm5, sximm8, status, datapath_out);
	input clk, loada, loadb, write, vsel, asel, bsel, loadc, loads;
	input [2:0] readnum, writenum;
	input [1:0] shift, ALUop;
	input [15:0] mdata, sximm5, sximm8;
	
module counter(clk, reset, loadpc, msel, C,);
        input clk, reset, loadpc, msel;
        input [15:0] C;
       
RAM #(16,8,"data.txt") RAMInstantiate(
                (~KEY[0])		inp
                (readAddress), 		inp
                (writeAddress)		inp
                (write), 		inp
                (B),    		inp       //B is what is being written in
                (mdata) 		out   

module instructionReg(clk, mdata, loadir, instruction);
        
        input clk, loadir;
        input [15:0] mdata;
        output [15:0] instruction;
        
        

//OUTPUTS ARE THINGS I HAVE TO WORK WITH
//INPUTS ARE THINGS I NEED TO PROVIDE

//GENERAL FORMAT
//first receive an instruction
//assign state things and next state things depending on which operaiton
//under each state, u shuld have another set of case statements describing what to do in each state
//after all the things are done in each state
//You should load the instruction register by enable loadir = 1 or something along the lines
//do this for all the operations
