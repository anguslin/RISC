module DFlipFlop(clk,in,out);
  parameter n=1;
  input clk;
  input [n-1:0] in;
  output [n-1:0] out;
  reg [n-1:0] out;

  //update on rising edge
  always @(posedge clk)
    out = in;
endmodule
