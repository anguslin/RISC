        
//module to display the value of datpath_out DE1-SoC

// One bit per segment on the DE1-SoC a HEX segment is illuminated depending on the input from datapath_out
//The HEX display bits are as follows:
          
//    0000
//   5    1
//   5    1
//    6666
//   4    2
//   4    2
//    3333
          
module HEXDisplay(inValue, display);
        input [3:0] inValue;
        output [6:0] display;
	reg [6:0] display;

        always @(*) begin
                case(inValue)
                        4'b0000: display = 7'b1000000; //0
                        4'b0001: display = 7'b1111001; //1
                        4'b0010: display = 7'b0100100; //2
                        4'b0011: display = 7'b0110000; //3
                        4'b0100: display = 7'b0011001; //4
                        4'b0101: display = 7'b0010010; //5
                        4'b0110: display = 7'b0000010; //6
                        4'b0111: display = 7'b1111000; //7
                        4'b1000: display = 7'b0000000; //8
                        4'b1001: display = 7'b0011000; //9
                        4'b1010: display = 7'b0001000; //10 = A
                        4'b1011: display = 7'b0000011; //11 = b
                        4'b1100: display = 7'b1000110; //12 = C
                        4'b1101: display = 7'b0100001; //13 = d
                        4'b1110: display = 7'b0000110; //14 = E
                        4'b1111: display = 7'b0001110; //15 = F
                endcase
        end
endmodule
